`timescale 1ns / 10ps
/* verilator coverage_off */

module tb_magnitude ();
    initial begin
        $finish;
    end
endmodule

/* verilator coverage_on */

